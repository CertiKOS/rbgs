(** Convenience re-exports for the refinement-based game semantics
    development so examples can depend on a single module name. *)

Require Export models.IntStrat.
Require Export models.EffectSignatures.
Require Export models.IntSpec.
Require Export models.LinCCAL.

